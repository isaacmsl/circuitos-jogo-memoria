PACKAGE our_pkg IS
    TYPE CARTAS_JOGO IS ARRAY (0 to 15) OF BIT_VECTOR(2 DOWNTO 0);
    TYPE CARTAS_DISPLAY IS ARRAY (0 to 15) OF BIT_VECTOR(6 DOWNTO 0);
END PACKAGE our_pkg;